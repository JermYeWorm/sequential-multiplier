`timescale 1ns / 1ps

module Sequential_Mult(

    );
endmodule
